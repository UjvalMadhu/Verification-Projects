////////////////////////////////////////////////////////////////////////////////////
///                        UVM Verification Project                             ////
///                           AMBA APB5 Protocol                                ////
////////////////////////////////////////////////////////////////////////////////////
///   APB5 Interface                                                            ////
///   Copyright 2025 Ujval Madhu, All rights reserved                           ////
////////////////////////////////////////////////////////////////////////////////////
//  CVS Log
//
//  Id: apb_inf.sv,v 1.0
//
//  $Date: 2025-01-11
//  $Revision: 1.0 $
//  $Author:  Ujval Madhu